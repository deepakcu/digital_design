// Design a circuit that accepts an n-bit
// grey code as input and produces the equivalent
// n-bit binary code
//
// Sample 3-bit grey to binary conversion
// grey  bin  
// 000   000
// 001   001
// 011   010
// 010   011
// 110   100
// 111   101
// 101   110
// 100   111
module grey_to_binary #(
   parameter WIDTH=3
) (
   input [WIDTH-1:0] grey
   output [WIDTH-1:0] binary
);


endmodule
